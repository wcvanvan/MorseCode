`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/11/27 18:50:48
// Design Name: 
// Module Name: converter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


// module converter(
//     input mode,
//     input clk
// );
//     // reg mode; // 绑定到开关12
//     decoder dec(.turn_on (~mode));
//     encoder enc(.turn_on (mode));
// endmodule

// `timescale 1ns / 1ps
// //////////////////////////////////////////////////////////////////////////////////
// // Company:
// // Engineer:
// //
// // Create Date: 2021/12/20 20:49:29
// // Design Name:
// // Module Name: encode
// // Project Name:
// // Target Devices:
// // Tool Versions:
// // Description:
// //
// // Dependencies:
// //
// // Revision:
// // Revision 0.01 - File Created
// // Additional Comments:
// //
// //////////////////////////////////////////////////////////////////////////////////


module encode(input clk,
              input rst,
              input [7:0] s1,
              input [7:0] s2,
              input [7:0] s3,
              input [7:0] s4,
              input [7:0] s5,
              input [7:0] s6,
              input [7:0] s7,
              input [7:0] s8,
              output wire beep,
              input [8:0] switches,
              input speed_adjust,
              input sound_begin);
    
    reg [143:0] code = 0;
    always @(s1) begin
        if (rst) begin
            code[139:126] = 0;
        end
        else begin
            case (s1)
                5'h10: code[143:126]   = 0;
                4'h0: code[143:126]    = 18'b0000_11011011011011;
                4'h1: code[139:126]    = 18'b0000_10110110110110;
                4'h2: code[139:126]    = 18'b0000_10101101101100;
                4'h3: code[139:126]    = 18'b0000_10101011011000;
                4'h4: code[139:126]    = 18'b0000_10101010110000;
                4'h5: code[139:126]    = 18'b0000_10101010100000;
                4'h6: code[139:126]    = 18'b0000_11010101010000;
                4'h7: code[139:126]    = 18'b0000_11011010101000;
                4'h8: code[139:126]    = 18'b0000_11011011010100;
                4'h9: code[139:126]    = 18'b0000_11011011011010;
                default: code[139:126] = 0;
            endcase
        end
    end
    always @(s2) begin
        if (rst) begin
            code[125:108] = 0;
        end
        else begin
            case (s2)
                5'h10: code[125:108]   = 0;
                4'h0: code[125:108]    = 18'b0000_11011011011011;
                4'h1: code[125:108]    = 18'b0000_10110110110110;
                4'h2: code[125:108]    = 18'b0000_10101101101100;
                4'h3: code[125:108]    = 18'b0000_10101011011000;
                4'h4: code[125:108]    = 18'b0000_10101010110000;
                4'h5: code[125:108]    = 18'b0000_10101010100000;
                4'h6: code[125:108]    = 18'b0000_11010101010000;
                4'h7: code[125:108]    = 18'b0000_11011010101000;
                4'h8: code[125:108]    = 18'b0000_11011011010100;
                4'h9: code[125:108]    = 18'b0000_11011011011010;
                default: code[125:108] = 0;
            endcase
        end
    end
    always @(s3) begin
        if (rst) begin
            code[107:90] = 0;
        end
        else begin
            case (s3)
                5'h10: code[107:90]   = 0;
                4'h0: code[107:90]    = 18'b0000_11011011011011;
                4'h1: code[107:90]    = 18'b0000_10110110110110;
                4'h2: code[107:90]    = 18'b0000_10101101101100;
                4'h3: code[107:90]    = 18'b0000_10101011011000;
                4'h4: code[107:90]    = 18'b0000_10101010110000;
                4'h5: code[107:90]    = 18'b0000_10101010100000;
                4'h6: code[107:90]    = 18'b0000_11010101010000;
                4'h7: code[107:90]    = 18'b0000_11011010101000;
                4'h8: code[107:90]    = 18'b0000_11011011010100;
                4'h9: code[107:90]    = 18'b0000_11011011011010;
                default: code[107:90] = 0;
            endcase
        end
    end
    always @(s4) begin
        if (rst) begin
            code[89:72] = 0;
        end
        else begin
            case (s4)
                5'h10: code[89:72]  = 0;
                4'h0: code[89:72]    = 18'b0000_11011011011011;
                4'h1: code[89:72]    = 18'b0000_10110110110110;
                4'h2: code[89:72]    = 18'b0000_10101101101100;
                4'h3: code[89:72]    = 18'b0000_10101011011000;
                4'h4: code[89:72]    = 18'b0000_10101010110000;
                4'h5: code[89:72]    = 18'b0000_10101010100000;
                4'h6: code[89:72]    = 18'b0000_11010101010000;
                4'h7: code[89:72]    = 18'b0000_11011010101000;
                4'h8: code[89:72]    = 18'b0000_11011011010100;
                4'h9: code[89:72]    = 18'b0000_11011011011010;
                default: code[89:72] = 0;
            endcase
        end
    end
    always @(s5) begin
        if (rst) begin
            code[71:54] = 0;
        end
        else begin
            case (s5)
                5'h10: code[71:54] = 0;
                4'h0: code[71:54]    = 18'b0000_11011011011011;
                4'h1: code[71:54]    = 18'b0000_10110110110110;
                4'h2: code[71:54]    = 18'b0000_10101101101100;
                4'h3: code[71:54]    = 18'b0000_10101011011000;
                4'h4: code[71:54]    = 18'b0000_10101010110000;
                4'h5: code[71:54]    = 18'b0000_10101010100000;
                4'h6: code[71:54]    = 18'b0000_11010101010000;
                4'h7: code[71:54]    = 18'b0000_11011010101000;
                4'h8: code[71:54]    = 18'b0000_11011011010100;
                4'h9: code[71:54]    = 18'b0000_11011011011010;
                default: code[71:54] = 0;
            endcase
        end
    end
    always @(s6) begin
        if (rst) begin
            code[53:36] = 0;
        end
        else begin
            case (s6)
                5'h10: code[53:36] = 0;
                4'h0: code[53:36]    = 18'b0000_11011011011011;
                4'h1: code[53:36]    = 18'b0000_10110110110110;
                4'h2: code[53:36]    = 18'b0000_10101101101100;
                4'h3: code[53:36]    = 18'b0000_10101011011000;
                4'h4: code[53:36]    = 18'b0000_10101010110000;
                4'h5: code[53:36]    = 18'b0000_10101010100000;
                4'h6: code[53:36]    = 18'b0000_11010101010000;
                4'h7: code[53:36]    = 18'b0000_11011010101000;
                4'h8: code[53:36]    = 18'b0000_11011011010100;
                4'h9: code[53:36]    = 18'b0000_11011011011010;
                default: code[53:36] = 0;
            endcase
        end
    end
    always @(s7) begin
        if (rst) begin
            code[35:18] = 0;
        end
        else begin
            case (s7)
                5'h10: code[35:18] = 0;
                4'h0: code[35:18]    = 18'b0000_11011011011011;
                4'h1: code[35:18]    = 18'b0000_10110110110110;
                4'h2: code[35:18]    = 18'b0000_10101101101100;
                4'h3: code[35:18]    = 18'b0000_10101011011000;
                4'h4: code[35:18]    = 18'b0000_10101010110000;
                4'h5: code[35:18]    = 18'b0000_10101010100000;
                4'h6: code[35:18]    = 18'b0000_11010101010000;
                4'h7: code[35:18]    = 18'b0000_11011010101000;
                4'h8: code[35:18]    = 18'b0000_11011011010100;
                4'h9: code[35:18]    = 18'b0000_11011011011010;
                default: code[35:18] = 0;
            endcase
        end
        
    end
    always @(s8) begin
        if (rst) begin
            code[17:0] = 0;
        end
        else begin
            case (s8)
                5'h10: code[17:0] = 0;
                4'h0: code[17:0]     = 18'b0000_11011011011011;
                4'h1: code[17:0]     = 18'b0000_10110110110110;
                4'h2: code[17:0]     = 18'b0000_10101101101100;
                4'h3: code[17:0]     = 18'b0000_10101011011000;
                4'h4: code[17:0]     = 18'b0000_10101010110000;
                4'h5: code[17:0]     = 18'b0000_10101010100000;
                4'h6: code[17:0]     = 18'b0000_11010101010000;
                4'h7: code[17:0]     = 18'b0000_11011010101000;
                4'h8: code[17:0]     = 18'b0000_11011011010100;
                4'h9: code[17:0]     = 18'b0000_11011011011010;
                default: code[17:0]  = 0;
            endcase
        end
    end
    buzzer b(.clk(clk), .rst(rst),.code(code), .beep(beep), .switches(switches), .speed_adjust(speed_adjust), .sound_begin(sound_begin));
    
endmodule
